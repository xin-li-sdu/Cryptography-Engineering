`timescale 1ns/100ps
module main_tb;

    reg			    clk		            ;
    reg			    reset_n	            ;
    reg             sm4_en              ;
    reg   [127: 0]  data_in             ;
    reg   [127: 0]  user_key_in         ;
    wire            ready_out           ;
    wire  [127: 0]  result_out          ;
	

    //always #1  clk = ~clk;
initial begin  
    clk = 0;  
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk;  
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk;  
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk;  
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk;  
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk;  
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk;  
#10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk;  
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk;  
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk;  
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk;  
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk;  
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk;  #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk;  
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk;  
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk;  
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk;  
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk;  
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk;  #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk;  
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk;  
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk;  
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk;  
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk;  
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk;  #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk;  
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk;  
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk;  
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk;  
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk;  
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk;  
#10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk;  
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk;  
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk;  
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk;  
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk;  
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk;  #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk;  
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk;  
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk;  
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk;  
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk;  
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk; 
    #10 clk = ~clk;  
  end  

	main uut(.CLK(clk), .RST_N(reset_n), .SM4_EN(sm4_en), .IN_DATA(data_in), .IN_KEY(user_key_in), .OUT_DATA(result_out), .OUT_READY(ready_out));
	
	initial begin
		clk = 0;
		reset_n = 1'b0;
		sm4_en = 1'b0;
		#10
		sm4_en = 1'b1;
		reset_n = 1'b1;
		data_in = 128'h 01_23_45_67_89_ab_cd_ef_fe_dc_ba_98_76_54_32_10;
		user_key_in = 128'h 01_23_45_67_89_ab_cd_ef_fe_dc_ba_98_76_54_32_10;
		#10
		reset_n = 1'b0;
		sm4_en = 1'b0;
		#10
		reset_n = 1'b1;
		sm4_en = 1'b1;
		data_in = 128'h 01_23_45_67_89_ab_cd_ef_fe_dc_ba_98_76_54_32_10;
		user_key_in = 128'h 01_23_45_67_89_ab_cd_ef_fe_dc_ba_98_76_54_32_10;
		#70 if (ready_out == 1'b1) $stop;
		
	end 


 initial begin
    $dumpfile("test.vcd");
    $dumpvars;
  end

endmodule
